LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE Constants IS
	CONSTANT VCC: std_logic := '1';
	CONSTANT GND: std_logic := '0';
END Constants;